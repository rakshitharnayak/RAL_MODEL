// N means how many packets to generate
`define N 2  
